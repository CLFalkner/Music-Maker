PK   �}�Sz���)  �    cirkitFile.json�ݎ�6��_eP{Wj0D�����Y{����M��P��va�U}�c<�t^�<�2����J��Ӄs���N�B��"��^�unv�ۻa���������#՗?uw�/��5�_�nv���/?]|���\=���P��ߦ6�vpa84]��UnT퍵�߻�>���������O�/߯@b�#1�T��j1�T�쬘A�`vN� U0�F� U0;/f�*�]3H�.��
f׊�
)F��X"Q B�<V�<X�%�<\�%�<`�%�<d�%�<h�%�<l�/�۟���7��p�>�j?Сr&�*{�:�9oZwt���^�<�%�<�%R�Lw��Bw���I���Zw��Bw��Bw��Bw��Bw��B;��B;�)���N�D���N�D���N�D� ����i�S,�(�S,�(�S,�(�S,�(�S,�(�S,avN;��B;��B;��B;��0@*��N;��B;��B;��B;��B;�f��c�X"Q�c�X"Q�c�X"Qؕ������c���L_E}ul��M��[�;#Ϣ�ٿ��2�Uw���v�ݗ������o���px���p�D� |咇�F���B���B���B��f��!\,�(�!\,�(�!<�(��&��9~��G�qD�����t&	BmGX�A�Kgv5�v5�vP:�ҙ����bm�����PO���vrX�;��3��hى��z.X�7X�C�(�{�]����f�X�C�Kgvk�����r�w���lĚ=b��#,�ٵX۵X�A�KǓ8�� 8���������ΤЩ8�"p2E�l
�G`>���8�����'+��N��|��i�`��s,��x�8�~�d�G`>���8a����'փ��<�|������F��8q!p��#0/� ăs,��x	�~���G`>^|��K�S8w���K�]�|��?`��s,��x��~���G`>^d�8w���������]�|��m`��s,��xI�~���G`>^L���?�|��e�`���,��x'�~���G`>^z
�z6z:8����Â�,��x�/�~���G`>^��8������X���?r����:��{Sy7$1��������p�뾎�x^(��x]9�����G|ﾕҩ���Xpփ�#0���ρ�,�����~��G`>.� �8������F���z�|��r`��Ӏ�,� ���`���%F��g=X>�qq���Y���|\�l?p��#0���`��ǥt��k�����|\l?p���#0�/��`��gN*A��?�|y���C_�*%48}i�����|\�
l?��~��~p�Ҁӗ��`��ǅ����/X>�qI3�������|\�l?p���#0����σ�,��� �~���G`>.��8}�����`��V����uu��C<V��56쇾s-WǱ����r:����nda�y�����J��ͭ����la�yA����J����%X��k�6�=-u��	�.������]�J�}/���������J��/ۥ���4�	�/�ӫ�����}�J��/ۻ��������J_\B���h*m/}�ڕ˦�V�a7Cz��ѩ��So�]X�N-|`��&���$�0�]�J���qg d� a! �|s�Ra���)m/|e{ꔶ��@B� �d{ފBɸ����-��~7�?���;�妴���,S�^��eۨ��>o��%��}�l������P�EGi{��e�b����������������/�/�/�/�/�/�/H����������������������#�B��B�k���
���_+��V���m\])K}�=(�,|�|X�RK>�ٵᬍ;����~l�[GF�܎���7τ�dm�u�����Nh� 3�ڀ�֑b���ߖ����,75_Wnj����:�"��Њb��E�EcD�=�΋�}�ė�'٥73/��̲q�e�%�|}�I�[�	��?�t�Wt�u����U���������ޘ���z�s�i��Umh��h����7~�}mB��g��|<�oc�����p{}{w��WɍLD�ˌ�\\J���x�"�����$d�ׄ!	�La�@B�;U"����$d���!	�b�@B�;�"�������ڸ����(%3�AL��M���R2cg����(%3NQ1�J�7�����	�QJf�Jb����QJf��b���qpX�aq�d��� &X�aq�d�i� &X�aq�d��� &X�aq�d�i�t�-,����8ĄI���⸅�q����`q���8JɌ+@L�8naq�d�� &Xw�8�R2�R
,�;XG)�q��	7&���q��(%3.Q1�⸃�q������`q���8JɌK`@�~`q���q���ꀘ`q�����g/���JƄF���(%3.S1��x��(%3.�1��x��(%3.�1�⸇�q������`q�����RyU�y4��XN
�J*���jv��hpU�]5XI����E��@�j��
���kA�U�v�`�֏,�I߱i��]神1�Y��
��y�g�*Ю�����΋Bc�:/���+���ݼX4\hW�l�_�E�1v����X@��TX�n^\�
��+���`��@'�R�%Z�۬c[��K)��ɻH'�"��K��thy���mu�/Zҡ�9�:����ThI������V'S�%Z^àc[�LL��thy-��mu�1Zҡ5'kߑ����Th� �\�t�2���ThI�����|X���ThI���*��V'/S�%Z^s�c[�/bJ��t�Z'/�u�2Zҡ�5p:����ThI������V'/S�%Z^��c[��L��thym��mu�2Zҡ�5�:����ThI��׺��V'/S�%Z^��31I'/S�%Z^{�c[��L��thy��mu�2Zҡ��:�U���4]Q'/�:y����ThI������V'/S�%Z�1�c[��L��thM����,Ҷ9-b�
�9�Fi[��L�6�K�����eV'/S�%Z���b[����В-�ѱ�N^�BK:�\EǶ:y�
-��rm���e*��C�5jtl���L'/S��Z;:����ThI��k��V'/S�%Z�}�c[��L��th����mu�2Zҡ�ZT:����ThI��kj�ض���ThI��k���V'/S�%Z�q�c[��L��th�V��mu�2ZZ���16:yY����В-��ӱ�R��2:yY���5:y�
-��r-C���e*��C�5ul����В-זԱ�N^�BK:�\#SŶ^'/S�%Z���c[��L��th�f��mu�Z�܏E�y�P�=�J��B��ڴ�*+�dK7����T�.TY��]��RݺPe�u��J�B���ϥ^r^���m�Z*��ߵ�UKe0���i�Ƈ׶	-��x��f��2����]*Ke0^��d�Ƌ�v\,��x�ھ��o]���X*�J�^�'�����5?���Z"3z����(�(�O����/���`�xmW��^�Y��o���Y��G���k����|�b��N�����;��ќ6�
��QvQ��~���E�u`b���Q�2/n0^���R�Ƌ�6.*���(ֶ*����MxJe0^���M�Ƌ=Ƌ=h|��������������������4̆��������������������-�xq�xq�����-Ƌ[��/n�zq\g����\�\���c�Um�m8�u_����z��I��%�T�s�.��8�}��t��������vΛ����h���+ڤRCXΎ�mRq��� �&���s���ȹI�l�ܤr6nn�:snXb��$�&S���&c� m���侧P��4瞃�����c�)����&����ћ�߷�(��]�B�Fv�}l鸯����\_u�>V��wvO~w~f�&�������9FW��M�Ma�j�|���&�Μg٤��Qf�p��������Ȗo��|7���]w���|G^��t�"���Z"��߀"��ߦ"����"����"��{"��{"��{2"���zE���ڸ����(%3u�0L��M���R2S�����(%3ML�0�b8��8J�LS�0L�8^��8J�L��0L��7���5,����4g���5,����4����5,����4����5,����4���⸅�q�����b�p#)��X��8�R2�`,�[XG)�ir2�	�-,����4m����QJf�Ѝa��q��(%3M5�0���q��8�`q�d��&Xw�8�R2�\,�;XG)�i��,�7�8�R2��,�7�8�R2����&��&,�7�8�R2�,�7�8�R2��,�{XG)�iQ�	�=,��)�׷��'�U�24 URa%V��j'�U�v�`%V���&�U�v�`%V��j٢U�v�`%֔w��5+c��+���~��]��h��
k꣨�5+_��+���]V��
��+���]V��
��+���]V��
��+���`��@'�R�%Z�۬c[��K)��ɻH'�"��K��thy���mu�/Zҡ�9�:����ThI������V'S�%Z^àc[�LL��thy-��mu�1Zҡ�5%:����ThI������V'+S�%Z^��aA'/S�%Z^��c[��L��thy͕�m���)}���j������ThI������V'/S�%Z^˧c[��L��thyM��mu�2Zҡ嵕:����ThI��׈��V'/S�%Z^�c[��L��thyͮ��$��L��thy�mu�2Zҡ�5�:����ThI��ׂ��Vi���tE�����eV'/S�%Z^��c[��L��th�ƀ�mu�2Zҡ�Z	:����ThI��k>��V'/S�%Z�]�c[��L��th���m�N^�BK:�\KDǶ:y�
-��rM���e*��C˵]tl����В-רѱ��J2��d:y���˜N^�BK:�\3HǶ:y�
-��r�#���e*��C�5�tl����В-עұ�N^�BK:�\SKŶ�N^�BK:�\LǶ:y�
-��r�3���e*��C˵�tl����В-לӱ�N^�BK:�\;OǶJU>��|��e�N^���e*��C˵ul����В-�dԱ�N^�BK:�\[RǶ:y�
-��r�L�z��L��th�֧�mu�2Zҡ嚥:����Thi��Vч�?���Uwp�r]���U�w����\��s��Jm�B��j��*+u�UV*o����.TY�n]��R��Pe��t��J��R�9/�{�6}-�����֪�2^���T��kۄ��`�xm3�RP�x��.��2/^��T��k;.��`�xm_�ҷ.Ƌ�v,�u%0^���^�Ƌ�6�+��x��q�2/^ۈ�T��k۝�ʀz�/^��T��k�m��`�xmO�Ҭ��k;G��`�xm�RPb��ⵍ�Je0^��=P�Ƌ�6�)��x��V7�2/�/���	�{�{�{��������0ƋƋƋ#Ƌ#Ƌ#Ƌ#Ƌ#Ƌ#Ƌ#Ƌ#h�����-Ƌ[��/n1^�b��=��up����np�sݾj�MW����X�}��_�6���O�T�ަ�p�>�d:T��P�`Ug;�M����W�I��mR�\�Y�ۤr��6����M*gC�&���s�����I�l���u ��x���l�d0�{�;�6����>��x���>�_�W�D_�>z������(�I��}�����㾢��+wp}���X���=�!�y�M*gY:כ�]Ն6�7FS���W��C�kBgγlRy���e�Ͽ�����������G[_^�ru7��\w���]��n������O/'-߰׈�;�/E''��Jx�Z���܊^�;�;����Sz��$���Z&Y/HZ��]�t2���)��6�����0�!)L���0c�0������/4����(��:���$?���$6=I���nG�'�ď���8ܐ$��,ԖO��|�+��.b18~}��l��E(�����:�K�W"�F+��N���݇���"�y�J	��W=���D�s%WN���)�¦����)"q�n����y��d%nl��+9��!���ҩ�:!Y�+���sE疼�\��[�\��[���Kߖ�IDy
$z��۠~��4N7�|����u7�Ҙ��D�������[�[A��W�(�A8�a�i��N�F�������'�~�'�7� ��J���7� ��J���7� ��J���7� ��x�*��E�|�o^�V���_i߼j�X��?�y�Z��w~�b�7�������Χ�^�!L�1��s1L�q�,�`�D��Y4�0�Ƽ����s�{��{���sn)�p:	�'��J0��%
��t�	�B:�C!�x�@�� ���P�D�&�Q�D�I)�7�� ���2��o 
�p�t�o2GN���#'���'+��
�I�;�xr��� ���#+���#+@0H��O��]
qB!�C(Ĺ	�B��A(�9�b���N���xʁ�S=�@��r��O9�t�'�m��@�٠ �P �tn($�O���|fib�H6{�����?t����?����v��ǫ��㯲���N��SM!�X��b	3VDR�%�XQIH!�0cE&!�X��b	3V�R�%�XQJH!�0cE*!�X�L��a=�?	@�f*�%� �PQ���ʂI9 q� �T�a����aN�!��T�V���v$�r �k�r3�$�@tO�S@x��U�a�m����Z«\�LKI9 ��W������r �i��r3m�%�,���\�L�{I9	?"��S��r3�P&� �S��r3�&� �S��r3��&� �S��r3�'� �S��r3�T'�@�"�P���\�L��I9 ���\�L��I9 ���\�LJG���S����<�r ��g�l�K�b�%��m�f��Q��� ��5̴���m@��k�i_K) �z@��k�igM) �z@��5�+`�z<�D�G`>�e���z�a�̗�TG�A��#0_V} ���/��<��aA 6��3�]=nV6�;�9�9�|�$����zx�9=؜X>�] �/����&�g�(����`sb��gv-�~-�~X>��Ht����		Mȓ9�6�g0���:�!t&$4!O�E��ɀ		M���6D�/`BB��e��9��Є<�mCt�&$4!OG����		MhNV:bl��P�����쳧��':g!t�&$4!/4@�y��0!�	y�چ�LHhB^���!����:m��iK�N[���&�5h��0!�	yQچ�LHhB^Є�!:m��c�m�N[���&�dh��0!�	yچ�<LHhB^���[��S���&�Ňh��0!�	y�$چ�<LHhB^�!|�|�:O��<Ţ�0!�	y�-چ�<LHhB^(��!:O��d�塂f������ǘ���w%����䄳{�@g1�ŀ		M����6t�,LHhB^�!:�����m��b���&�Rh��0!�	�Lچ�5.�,L�%.�6Dg1`BBry��Y��Є\ZmCt&$4!�EA����		M�%]�6D�)`BBr9�t�&$4!��A����		M�e��6D�)`BB��>16D�)`�|Sӷ�-��败A�-`BBr�(�������iK�N[t�&$4!��B����		M����6D�-`BBrm4��i��Є\�lC�N[���&�th��0!�	��چ�%'���-N�.��3��X�>��X�>�tX�y��}V���}Va��}V��}VѴ�}V���}VA���(��|��R��{��
H�0��T@���c�RO̷�*�B�'�a�
H=1��T@���O�RO��X*}�I=1�ըT@�Z�Y7�H������o�nT+ѓ��]�Rt�R/�w�)�Y�3=�R=��|�-bJ�}Oi��wS)��c%y\��&J�b�$zm��z�6!��H�o�Q* ��|��R���K�
H�����h�o�P* ��|ӂR�'z�'zq6/�D/�D/�D/�� �� �� �� �� �� �� X�zb�zb�zb�zb�zb�zb�zb�zb�zb�zb�qJ=1J=��zb+��Vꉭ�[�'�oxb\g����\�\���c�Um�m8�u_�n����$���ѕ\g�\�yDb8�6و�31T1�C���yӺ�3v�bO�P)��/�tK�B��b�J.�In�h�&���&'��ǚ�Ʈ6ɽO7�#�nj�F4����`��\{%�ߦ���+qa�ނs��mz�-���7�B��X�Jl�i�x<V�Q���h���M�i�}K~)L�<}�����ӷ��cK�}EG_W�������:���{�C8��>�oj�Ƌ�s�i��Umh��c4Uk�}�?ľ6!t��oj?���ˋ�vW���v��/>�z��]|�����f��l��a�Q�Ǉ]��t���!���qx���m������9��jnQ��ܢ�5���E�-jnQs��[Xna��q����[Xna����[8nḅ�n�nḅ��[8n�E�-n�p��[4�Es��[4ܢ�����s�-<���v��[xn�E��[n�E��[�Ѵ�"p��-"���"r��-"���"r�8�n�E�-Zn�r��[��"��>�e��UNoj�%N�|&�n�s�r��`˓y�`ˣ��Az����fx��h�~L2��Ss���4�ϊ�D�峨r�fo�[@�m.�q'4��[�́��f@�"9aX���7ݼ�KN%t�gs^(�k%t�Ϥ��i�Y�٘��lu�F��T ��gs�>��W�ƬY������`c.�.��8	�h�l��n�e�q@@4&��"�_I��~Q�q���t\4a �Y��[�y�|�g-�oM���,F�oXC�:��x#{�����?}�]w�ᚻ�3h��������~�O������&��=������o>�-<�����o1��}���~�W������f�OOVɍb�����<]w~���\��̓Er��'���0O���a�̑[���A�9����,�����Cuus��]_�?��orI����?�=�I�pr���B���a�p�O�� ���{�1�_ǿ����/����0������_2�����͏�D7���g����/��#���uo��E����n���?'݋����~H?�w�uu�����n�ߏWwC��!a'3���<�����p����^����W7� ���:~WW���jKj
�į�k/�������ɲ��I�b���VƦ�|?����PW�R3�G�q8������9Lm6��]^��]�[�M`��/|'Ww�������2�ړ>_~�u�n������a�:>�$p�D.f����z�8
ێ�O�ڄ��*�y���+zU=�Gή����$��0q�`��8�`\64���{S�5�x�=�S�k��L8{��E�S۞�o��qN�x\�c����x����/��|�e[-fc�-�	�q�ͩ��曙+�	�;9��E����=1iXVˏZ��NNJ�i���ܩV�|T�E[��vW7i�M�8>����5�����:��߄�&;��'��9T�D�E����a�m�8{�W���E_�����Le尹E�OV��m�B��O[�h�>+�pQpX��[fEa�a�I��a�%A��J��-	ֳ3������̴"�x܂`;;�]֛�v���$7?lM�o���W���(Ͳ���5<{z�������t�m{��p��Ş��"W�9ɰ��˂+.I��F���$���+O��qK�M�Mp�8���B;]��}}
�h��0�|X��:2)ê]��T[<,Wk�I_?w�����nJ�������ǔ���᱿�����~������Ҕ������K4� Iy����<''�>���䢓�/C��<=ߋ���w�oҝ���XW����}5=�&�k�yJ�iŦ���W�}��S���9��n���4N5�֞�]�����7�#�I�v��|���u[��O����>$_p��i�8��=V�f�U8R]��j��;�D�q���E6͘�����A*ۼxHe����oG���|L����S��Cݾ�O_<���<sy��YS�����i�A��sڤ�O�P;��m(�5��2 �0ϒ�~�Y��yЂ���;<i�sO,6!>ߕ�z��}}e�맭w}��6=9�����`�>ݩ@��M7Y��i�4alS@��Q v˃L��`ۧ���w���W�{��>���ѫ���Pm������gvG��s�-����n~L�?��6u�ҋ�n\rl�Ԥ������nN�����+��Q/������~� ���*]����O�����?��g�����w����w7���|�c_Q�@��إ�t���Ylp�4�F��uC}M���f�leܐzM�T٣s�M7w�MS�{w��O��.��rp�]:������n����};�v�K�|�X��&�ns�E��`��[��87BJ��9G���� PK
   �}�Sz���)  �                  cirkitFile.jsonPK      =   �)    